////-------------------------------------------------------------------------
////    Ball.sv                                                            --
////    Viral Mehta                                                        --
////    Spring 2005                                                        --
////                                                                       --
////    Modified by Stephen Kempf 03-01-2006                               --
////                              03-12-2007                               --
////    Translated by Joe Meng    07-07-2013                               --
////    Modified by Po-Han Huang  12-08-2017                               --
////    Spring 2018 Distribution                                           --
////                                                                       --
////    For use with ECE 385 Lab 8                                         --
////    UIUC ECE Department                                                --
////-------------------------------------------------------------------------
//module  mouseclick ( input         Clk,                // 50 MHz clock
//                             Reset,              // Active-high reset signal
//                             frame_clk,          // The clock indicating a new frame (~60Hz)
//               input [9:0]   DrawX, DrawY,       // Current pixel coordinates
//					input logic [9:0] XMOV_MOUSE,YMOV_MOUSE,
//               output logic  is_mouse             // Whether current pixel belongs to ball or background
//              );
//
//	 logic frame_clk_delayed, frame_clk_rising_edge;
//	 logic [9:0] XMOTION,YMOTION;
//
//    always_ff @ (posedge Clk) begin
//        frame_clk_delayed <= frame_clk;
//        frame_clk_rising_edge <= (frame_clk == 1'b1) && (frame_clk_delayed == 1'b0);
//    end
//	always_comb
//	begin
//	XMOTION=10'd0;
//	YMOTION=10'd0;
//	if(frame_clk_rising_edge)
//		XMOTION=XMOV_MOUSE;
//		YMOTION=YMOV_MOUSE;
//	end
//    parameter [9:0] Ball_Size = 10'd4;
//    int DistX, DistY, Size;
//    assign DistX = DrawX - XMOTION;
//    assign DistY = DrawY - 10'd480 + YMOTION;
//    assign Size = Ball_Size;
//	 always_comb
//	 begin
//        if ( ( DistX*DistX + DistY*DistY) <= (Size*Size) )
//            is_mouse = 1'b1;
//        else
//            is_mouse = 1'b0;
//	 end
//
//endmodule

module  mouseclick (input         Clk,                // 50 MHz clock
                      Reset,              // Active-high reset signal
                      frame_clk,          // The clock indicating a new frame (~60Hz)
                      input [9:0]   DrawX, DrawY,       // Current pixel coordinates
                      input logic [9:0] XMOV_MOUSE,YMOV_MOUSE, //position of our mouse
                      //					input logic STOREBEGIN,STOREEND,
                      //					input logic [7:0] X_CHANGE,Y_CHANGE,
                      output logic  is_mouse,          // Whether current pixel belongs to ball or background
                      output logic  [9:0] Ball_X_OUT,Ball_Y_OUT
                     );

  parameter [9:0] Ball_X_Center = 10'd320;  // Center position on the X axis
  parameter [9:0] Ball_Y_Center = 10'd240;  // Center position on the Y axis
  parameter [9:0] Ball_X_Min = 10'd0;       // Leftmost point on the X axis
  parameter [9:0] Ball_X_Max = 10'd639;     // Rightmost point on the X axis
  parameter [9:0] Ball_Y_Min = 10'd0;       // Topmost point on the Y axis
  parameter [9:0] Ball_Y_Max = 10'd479;     // Bottommost point on the Y axis
  parameter [9:0] Ball_X_Step = 10'd1;      // Step size on the X axis
  parameter [9:0] Ball_Y_Step = 10'd1;      // Step size on the Y axis
  parameter [9:0] Ball_Size = 10'd3;        // Ball size

  logic [9:0] Ball_X_Pos, Ball_X_Motion, Ball_Y_Pos, Ball_Y_Motion;
  logic [9:0] Ball_X_Pos_in, Ball_X_Motion_in, Ball_Y_Pos_in, Ball_Y_Motion_in;
  logic [7:0] w,a,s,d,space;



  assign Ball_X_OUT=Ball_X_Pos;
  assign Ball_Y_OUT=Ball_Y_Pos;

  //////// Do not modify the always_ff blocks. ////////
  // Detect rising edge of frame_clk
  logic frame_clk_delayed, frame_clk_rising_edge;
  always_ff @ (posedge Clk)
  begin
    frame_clk_delayed <= frame_clk;
    frame_clk_rising_edge <= (frame_clk == 1'b1) && (frame_clk_delayed == 1'b0);
  end

  always_ff @ (posedge Clk)
  begin
    if (Reset)
    begin
      Ball_X_Pos <= Ball_X_Center;
      Ball_Y_Pos <= Ball_Y_Center;
      //				Ball_X_Pos <= {2{1'b0},start_pos};
      //				Ball_Y_Pos <= {2{1'b0},start_pos};
      //				Ball_X_Motion <= 10'd0;
      //            Ball_Y_Motion <= 10'd0;

    end
    else
    begin
      Ball_X_Pos <= Ball_X_Pos_in;
      Ball_Y_Pos <= Ball_Y_Pos_in;
      //            Ball_X_Motion <= Ball_X_Motion_in;
      //            Ball_Y_Motion <= Ball_Y_Motion_in;
    end
  end
  //////// Do not modify the always_ff blocks. ////////

  // You need to modify always_comb block.
  always_comb
  begin
    // By default, keep Motion and position unchanged
    Ball_X_Pos_in = Ball_X_Pos;
    Ball_Y_Pos_in = Ball_Y_Pos;
    //        Ball_X_Motion_in = Ball_X_Motion;
    //        Ball_Y_Motion_in = Ball_Y_Motion;

    // Update position and Motion only at rising edge of frame clock
    if (frame_clk_rising_edge)
    begin
      // Be careful when using comparators with "logic" datatype because compiler treats
      //   both sides of the operator as UNSIGNED numbers.
      // e.g. Ball_Y_Pos - Ball_Size <= Ball_Y_Min
      // If Ball_Y_Pos is 0, then Ball_Y_Pos - Ball_Size will not be -4, but rather a large positive number.
      // Pay attention to the velocity. We must always make sure that the ball only has velocity in one direction.
      Ball_X_Pos_in=XMOV_MOUSE;
      Ball_Y_Pos_in=YMOV_MOUSE;
      //				if(X_CHANGE!=0 && Y_CHANGE!=0)
      //				begin
      //				Ball_X_Motion_in=X_CHANGE;
      //				Ball_Y_Motion_in=Y_CHANGE;
      //				end
      //				else
      //				begin
      //				Ball_X_Motion_in=10'd0;
      //				Ball_X_Motion_in=10'd0;
      //				end



      //            Ball_X_Pos_in = Ball_X_Pos + Ball_X_Motion;
      //            Ball_Y_Pos_in = Ball_Y_Pos + Ball_Y_Motion;
    end

    /**************************************************************************************
        ATTENTION! Please answer the following quesiton in your lab report! Points will be allocated for the answers!
        Hidden Question #2/2:
           Notice that Ball_Y_Pos is updated using Ball_Y_Motion. 
          Will the new value of Ball_Y_Motion be used when Ball_Y_Pos is updated, or the old? 
          What is the difference between writing
            "Ball_Y_Pos_in = Ball_Y_Pos + Ball_Y_Motion;" and 
            "Ball_Y_Pos_in = Ball_Y_Pos + Ball_Y_Motion_in;"?
          How will this impact behavior of the ball during a bounce, and how might that interact with a response to a keypress?
          Give an answer in your Post-Lab.
    Answer:1. It has been updated when Ball_Y_Pos is updated. 2. For the design "Ball_Y_Pos_in = Ball_Y_Pos + Ball_Y_Motion;" ,
    The frame will create one delay so that the ball will go through the boundary for a while and then back to the screen; for the design "Ball_Y_Pos_in = Ball_Y_Pos + Ball_Y_Motion_in;",
    The ball will response the keyboard immediately and there will be no frame delay for the ball moving.
    **************************************************************************************/
  end

  // Compute whether the pixel corresponds to ball or background
  /* Since the multiplicants are required to be signed, we have to first cast them
     from logic to int (signed by default) before they are multiplied. */
  int DistX, DistY, Size;
  assign DistX = DrawX - Ball_X_Pos;
  assign DistY = DrawY - Ball_Y_Pos;
  assign Size = Ball_Size;
  always_comb
  begin
    if ( ( DistX*DistX + DistY*DistY) <= (Size*Size) )
      is_mouse = 1'b1;
    else
      is_mouse = 1'b0;
    /* The ball's (pixelated) circle is generated using the standard circle formula.  Note that while
       the single line is quite powerful descriptively, it causes the synthesis tool to use up three
       of the 12 available multipliers on the chip! */
  end

endmodule
